version https://git-lfs.github.com/spec/v1
oid sha256:dd48865d889d9b91e5e0aa94d40806df16591ab63b294b89108f9d5d7ca98eb4
size 2602

version https://git-lfs.github.com/spec/v1
oid sha256:e5f3fc806899d76a0a6e723478e1a07198546451f8258d3d660f8fa1fa319a3b
size 4631
